`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 1000
`define LAT_MIN 100
`endif

module pseudo_DRAM_inst#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/DRAM_inst.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency, 
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:4*64*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 1, DRAM_W_LAT =1, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8191];   // addr from 00000000 to 0001FFF


//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
Gj5FWUoMEla+h9opOdl/8JxGbAnYVz8uAGpppX6LBvYwxieoWLCavIiUDyyq6Gh4
BU7p02rY3qmGQECGXoDU23x54iSJDEB8MQZHX5dJs+nplLK1FQ5JpHWR37g9Q77x
XL2MRTppHDNSZXzTWRtSpFyyLi28cwIWXlO8jFuIgW0vgYGE2uvot3T2NA++eP9v
MZYugUIhEnn1/vQhnWBqBKif/x6YGFNnpXsBEzDprHhiXNvR1NWaFhubBISY2uAG
iR6EG9p969YMW02qy7DfilmzBf6hMTBNKU/leZW73k9TlKztM5DzHBLraGQrAClA
+t7gaPNkHrxmYjV5TOmuXQ==
//pragma protect end_key_block
//pragma protect digest_block
m/5G7OjZ+YuchIs8GdLy0NEv52k=
//pragma protect end_digest_block
//pragma protect data_block
4MWFx0pcYpj3HKdjpbThXdAKIvsUDPAfxA4vPEL24D5bD/rUe+I8Dg7yTay7b2Y7
CsiOzIWRU3LC9Vo28xQd6O0KVrXLKiwyff3JwtsJ0rS/KBQZlnf2lTHUgrSSrsgr
9k/Z5kC0qjRhlzGken1nLSQB1bRSFvr3XVIBslB8uzUmvvmUvU7vmcsZmMImsqDr
Qo1PD27qrkfIz7RxtSVZUtTAJvNiBbJlotrcw9gsu3kdji7dFyqJ5CTiHDkrdx9+
wLqyReAPxnUlN6sSVR5qjPgLONuJe2x5zAcOrNfIeA1sB1rJMhjjaOKXafF5zVW/
JWKHIngKVPajDijy2lCngpFMJZS7mmSLWDEqbXHqpBLvAFPVSn4Go/eoxPZuhg51
Nif9PP3jux1D7mUNQnV3jYHY6bw1kKarUT3rCUXwRfKENSuM00JsJMwTFfTD/rE6
6gtXxm3qu72+fdv7avV8nLG5hJrUoYBMLeDseL2iMiQOIKg+DmQa2wWj5dI0sznU
07dRNyJmGfmmPaGF6hvkkHlHmXfoSac3i4Od579kWs00cBVt4Ki5RLNcerbUn0AZ
jeLFRoPlAgknIGdBvBWu6I/doDccHQignm8caawwDZzcZyrCUWP89C+36Lpku177
RKomxWb0ciHdKsmuOE486EyU7JGkqSPvfmmlwyI4VB/8NnJpUxN3e39SnVKxZ8Ih
9PEL1fqrKFjM6/jrsDcwZ8Qx5AzOkPUDZ+RexL2wRiOTG20sGdpQ+6qJ74QfwXVC
4dkBYzyD/LKKI0Q4JZ4eRXz0ZXxYNcMQEp4eeEl4hSRb0U7gZtfirNpaAVodufIv
/+U//hAcWKUQVO20oFLZav6deBMgssYeeL6Lwdpaepgl//xWrxOrBA5muNMK7eJd
Q07JuaB6yVMB9UQX51C8aJsvbJ8n9B/DAKF4MpTpt4nFBBN0giRG8P7njByXpdcx
06649n00wPsTx+bgZqjJ9g8ELgMD0pRJqjw/HqZ/w/b3Vs7xPOo4iSDQxaBr41z3
eDHlgy82XfiAyFV7splTiIsfbfGh4y0QWfHB2TbfVIhED0yyIEuCJYA7FU2d9rL7
/urJXDNaBWZH4/RgQXQEvkwTpv84ZM/eSjyJ27DBrvQHF0TtPDvZ9IlTPcH9zwC/
KJNDawHJq4iegI7uXLpw9tlCJEadWgVeEW+0XCC4ippe8AoHljOrawmZJEEXMpz8
UN/4KlyN4fKI4ePU7PGnT2ZlQ5+FoZrAd6T3IlfPVPIBxLEuh94C/FNHho0alL21
1+BsDXCv/7N+LBrUMgzjHw8qMzX1PUZ996847Jyb/xdp4PpIpO6pAe/+gigzoii5
ZtS+BWZ8uzV/5ij+1f4CvqVmGQT+iHGkroOAk8I9SIMZ0G9f3q2KMy7AgUh8z2qJ
7B45Us1RMLyu2ltZXwenJStn/eUAlzGnUTb7k5Ok/5TGjAJn1zFuvYB6eEYy/3/J
Zz8Two7L1ulBdLjGgghHedSCOmPQoNVve9rQwfb5GUY9XHqBvFdu2OHcD4QXrw/Z
1LL54tBn9lzS95gMNVO0W89P/nB/Kf7OLObCfZ6S8vg5OYPaCqHR8L+5WJ2qYuCV
8lxwWuEFLEk27II1h2rVuCPSEt1i5rKcL6MkwaukQijOZLeayYzeCEj2Y69Ios40
X3UHDI2slt6DyMilSMBcLuQOWnSRtTLJFi2z4XR7X+bzNwJ+Mb1O9iVKn1735SFs
33kvclUHGxF6mRe9YOpaQQbBgL3vRkaE++mRO5RRIk5j9h+WBxKKj1YEYVbe7NsZ
cNzF44Q6ThR4e+7AVdDaqVFhPsbFaKohONpTkWC8kZNoptkFZm0FcPEEzh5nYv/v
gGQMbshF5FyWNiktFpj1OMpu9fvxCiWM9n7Jtx+HdfFuRtbWY+ErJX9qVh3sqIMI
wsW2hwh5r7xJEf4MlydKM9jF29zMYSME47hd2uWQ0ZzE3p0F9jX5tEU9yP/qQciF
H70heod+soLMwPl5D+Zl0Wl4WLa8vJIR989Dn0gxbbe73e6rTh19MIDg/R5tkpVa
Y6dDZ7JDGPV6W7MeQQLNUJiAXV6lhDjbv92Ccz96amxLUtqqITNqivZrNN3H1H3Q
5tZJoUqeve4jalOsJ486vzsZuCRMcyN0qkD6zqkxdnSAnyCUKAYs98/GdqMIuMhj
oNRxhMQZts307/RAhDWruVxsvL4tdelYsVrtDFZfu/RmPvilQ7JsojwKaRGVxH9B
pRnzsjB9lZWIeAm7F2KdLAeg2vqn+zJJPdG2ni92BgF7BOEfd8PutO8aTUUsbl90
Q0kRu3RFEroz9jcKiektLz3QP/T0TQGzFvTDQXO7q4C3kzmug6XLCs0Np6vzyGLG
s8LTqo020gHsUXvS8jJnl0dXshVuiCfUNdA+9dmTgueGtVeP5Qqir63pAok+SKm7
ap9WqTAl8GB5D7zPoR5THM+jLKRCJQ2JJ3zEMNLfA7Z1v/oGhy2peVGTuJMShw1I
BJ0ZUfPZC+7sgyS/42901HxQv3Q8HQVef2RHEhH9Fz7Y6gYojViV/9FQtojKqnyv
Grz9vCJRb8NLSQA2nsMC6l5SmGJGMBdjEmKNRLzgkEVM4VVesrG2zHaww2u3+l/6
IXzaM2nm3shFfZu8S4ZjKeG0/fHWEWdfpX1DlmQbKJZsCyFgpt45KHpzvun8+zsV
Zulbg4niN+i5w/W6gyywUU47BtXDdiQMm9590xwzeJTvMqjt7C/u3+CfAeHl7DZp
JDFlaAo1lFOfRH3EZg+qprndVs5cMjLG0ywsvuJK9G2In+v0xxlcJ5JV467gpSXk
Ujng49U8ZY+VrSO2KMAovc04dS/nDeNy3iUdNBLiRfmjBzeorIyk8Rv07YOgWVrK
RwZ2VSQDV1jN7JF3iQxnRVpOjWBywtrbPDrjYIPdgvw1/e0iWdF6uaQhG0SPKxo0
FLrICN09smwTK2CMbw4+qqpqfLN8vdfbZCX/AGij9xDjvm0Ok6u9aTpydCvSICn6
Wom2H9vFsiDf5Z8dBjibyT9bIF3mGtT3WMOhuReTEufXprfWOxzzVYnfmc103mYp
fAR69o2jq62rgDUmnK2de+HkED39spWgGk8Edzk6cItYWbGQaumLTp86yZidCQxy
duxJUN6ADCybY5LCS88mLh+aHjb4ZMtSIL7jhUpwjB4mhM4jJFFlZ2pNQ2UyrnGR
d8tEn9UfSb1rHxXOnUfFn7GnvbRiSF1b6LJxM6Kmy2ksh7lVwmlhk/pQI5Nspp9m
Fcwmf1p1CoQOVynFQuwAhyRxCWrRPQBBgBj7XnM0SftZ5PfzGoTqCk+G6onSccNK
UupFGWGmveoTjSRHrLIwSFKq8Xjr3B+JEp9ykvV5oWVu4BDrbvk3bsYv5svAnro6
lU3LbeC4rO+16ewjKbFhXqre0P1ZwQjiOmk95JIUcj9KVq3yGXKiJuXt5ZJ50cdI
SI6ShQWuBztXS1iVPgWvNrRnWgBKOTA+bZXLkBEQBkx3tSi1Fb5en9UahArI+90v
O43yORGxdKmTAB4o0heROgTwkki9K52KqPOGDLvBTDfDpgzezFBdXggTKVx2L8l6
fFU2Y8tM9LYhv85/nkOfubUlZ0HoODEgVw4Ny8JS3cYDeJOBRnCO9Ecm+K9jxOTQ
yFdhXEsPE60mC/WDm1GNptSTvGPNWfjFnZAwXLZIJX4DYH3sRkQvB9t0FBQi7diL
n44oCHKhdsihgpNm1v6N235MEopuU7yx8DOuu/uJxTUHVexNum1IA2e8rsf6EElp
l8W1Dmui/E+2/ZHFNv8NN7dRoKwHaUDpsJKqbmgOOROZDKd8ofVTb0aFtdQJbBPl
znrEUj/ZESwGoZI1B0jZktVBcrqn50ywgfcXekh5ymWgoQPbKO/2fnqp74uAqZzY
6EwcrIi3TRnEF078xHngdjer2WHcMe0R1LmqXpmhHwiHxcZp4B7kQDE/4ICbKojZ
kf9oH1S1IuT+hq7e/xjWJGPImGYuqboB4JIRRYwbkrhegK6JTj7wb1x3w4dZDnrt
lGNwDAZafSNDJAKu0HWO1qWvoc5khvKYpOxkULFVzR2BJa9+wbEX3nc69FtWtPqv
sdybUgyqT+Io4VfTJFYt/lJkeqqp6j5BbNLgmyg1Sbch3pZ1pBORNzS7qqNHR3nm
9pu6Qhq7s8cga5E6FrYRVJqX7J00KdshkRJvnMbqtqzPqShl1HYvXmsvztujHP3t
8WhU3k3qXzEA8GgnqBxF6wd8dqHhuw4EHGjxBeihpyw/C2Bh4tWIRiI9dENEA/wo
7ETfwxMzbcQ+ThDI0eglO1wvVrpKG2R2YQvbjZIUXiG90MIOpFJt5BluEmiLFRmX
wwYEQHSN1+D1kmaA0CgyBzA7NQf4G3WXKc9uu6dOfGv9bqlGpJ2mWArmsAWnVne5
sawJQhuIqvGpgcxK8M5zQMh4W8TKAkJfQ9lbtgL9f0bvfL+bZumCwSPuy12F+mw9
3KqOqorMgGBAGMO8W+blbHp1CuMgORSMBNi4q9hKp2b3kzYC6iTBAjTLtffGE5n+
yX0uOSyk0xsK4A8+VXNz/NfuMrlD9wTbDQgfkG3rnPCV3ZCe9cVIKwYqYBL4owJR
Nzwi9bYPEFLv0rNgFs/QYUOyecwBvyPF9ZVM3KPyRE6id+tvhXJZMuZQ7bCWi+A/
skJqAz+xVk9zjSlTrO9sNvyB+pKefphdskopcttsbJfv51qyo+O07lbg7hWl7UBy
yf4jnHJrJt37bug2gPfC1cT54LDNryRH/5VKEgXbLx3TZ7hvYROVEWkLyqk+izTb
cOCfZJGoZYIAf2hiSkPx4j81X2wY4OQQVO7Ds0tF62OMOyPSuYj2+/Rh+p1wgF0C
w7EaLNj4TTda6D4ROHyHzyL+TvMM1A3SPqsmJdXQJiBmrcQUfErj4gdsf6E5GRhW
3Jh9/LFBIWxI4mf0wrIwq2YzEnlbcN3JUgAKrOifefpb78YrzTxvjripiEAKA4mM
RHjg0X+txUWRj5f+q2QqZO/IuL+RXmEswfZCxKjL7AMtPKKBHdX03iz9WBXMwyKb
J+FKHTTwrNMPGgb88u0IEehpIp9qfjdxIPw/zFqrsSEWDHoV3tHsEzTMR4ujvWjd
WrerrLclevg0EWc+ljMhZpK/tEmby2EeOk3hb8JBY3dDydIUmtxUAxz1lJjXZmPu
3yC0n97+/JyCdBdcpdSNhNMBx96iN4CuhdVCqnMkKjgjd2ud/ZuBRHDdftQjNYuS
9J8eFzLLqi/vNX/vtO4I1i6ujKx0dbuJW2CqYAHiWQFLd/Iv1jtC12iMmzVemxDs
2JKj4C+N2QpCs88b2XpFLImBZt51220uJd+Vsxi3EETxTGAXNSV/SUKajINBTHLc
Txjh9PW2fjKAMLA6S4Qm5YD047+K2fEIsNpREV2jes2Ik53XZw+KleIj5geo/lis
ARlbbzO77e5OLSn2CO2hDf9VMdDTROl8U6K/x2wt+YtLxYdQvnR79XPVijGLdvWI
IrPqZ2LL+D4Xav+lofcdoZuyiesjiShmxC+L0opuGHArH1V9c+plB4tEpF6uqeew
AaOFQBgsBQ1IIUsZNwxWNNo1OL26Lt1yrFxr6rrq0H+EICdgm1lbYqH0EiXqF2i8
7Ch/eASGoht4cVDQUP792m5wusG6QX9a7EVI6zVwdtNcjTACz88rM8NVvWyUs31V
K6qw6YeIvpeuCLwGjzamuqp09Ej+CkNfXjjxEqIMDzvjCK1k2XmrzemfdFoWDK+S
m3LUJR+eu+tVALfmFBT6DGvqV2ljNvFv8qoVFhyW8NTFN2ZFu7sJpT/G3SpEEZMx
ua2RZ0ck6ApYaMFflGMgHUPC3UlLI5XtlhlaTU0aO1l2GrbO0HmqDK6vM2ViIwqn
8Affi2+CxiIikc0ahWg66bTw8oWwTWyUjn+N38ROu19O3WiFR65IaCXYsubc/hlW
WpCJN4LY00w8nAbZJ0H6ES+b+BtMi1ymw6WL7gOwxg77c0kvs5Q0R0GK472/2Lgo
7yJUqVojLEUTyG6/X1aMIf/avlFFu7vJVjPHFdAQlfRUEmhLqLYoYPXKK3z/cr9u
6fKnovQMgGyf3jILjHiT7K4QADWBVZ9nCSa+4wi8r+/qlDm9cxndjuHU0f26jvKP
5nymzRzwBalxfIxavT3eGsYG53S3z5X2TzvSxoNwjHN1UT7tQV0DLPixhsfIHVj3
BEiYL/uNAhPs1gMl5AkOgcyonusMrbt4tKCsJkYHX4FkXsXuNnYJLuDS0yO6lZj4
2CTVL8+zjfH383Zrlk9eVGTTsvbdh+0pPDnWqO96jloCEv0XeEw7Odw2WPnygrMq
ptYlsnvoxNLpgFW9gXv+yGZMspVrhyc6ah/Z6SpDr9MuPVx7Y5rP4vJxb+A3DC7n
ViDUjU0eNIK5YFK2PnQq4SyyQRKp6B50P7UBiN3jngXjg2IMPhnw3v6LYofRVbSV
S+TreVblZf3wePvGuG51kr1Rp+S783wG/SQei0JSD6nERezzqwBfzj6d7OsaJmAW
AmGq6oSFdkWxh3xYl1WhQb8fnOnpQ29adyWrYrSRobqkWMDLkSFV54tFeUfdovtD
wyt9ah4fednvaMrZy2uyzGNdRbgghD5w4RO2N+L6mBgGrCwO4D3EsqEJOl49tiTY
AILwT9kbpLZ1ggztC/I4pSmR+1SoroSQJwOyuPwYU6YQeZTPSUrsDcyHP9lTpyzd
TInfh/9cEKjTDV8I1sZ+aPTQD1nbeFh1sQNjSKz7uTr0bDcSLG81ISwPFtTxiRe7
2BXqhVECevDbrkSKaWv4pdoxcS1TGfrD5+uG5rQzQIBb1H6dKWwfyacx5l5tKQU9
o/2iFvbH1ifjr+betXAKN97LXgvDnN1k7YA8n5tm8g1SphoVi4EsqOYczejKuzP1
KMNAQW8yqGDeobd21xbRAySG1zZVx5peb94goz07aRs7fapyyEU2Dtx+qvvwAZbj
T55xAvx3Eo2ywQaPibSCd2T7+T/6WHPa2ZL96ojzBMfm5ygYpuuTYVPEEe4hjRP/
sFJuH0PC158FgfNEAR47fPe48kZFIArYYf+yw0R/o9Dg6113X1OxbnMEf16U0fXs
mAxIVQLAv3mKiVIPCxjV4mTIcryYyYZPnJf3lBrnzx6nHTt8rnXlH0FDJ9ckJOu4
j3VpiiiXY4IIxcsyANrL1uTXMsvRZWvxw3aiXqQ6Jf8Q2azzwWQfucNUOEngrA0M
bUk6WhMeRX2vGGU+2cjjSzj/klLRmyPf8U2oK2hPM5gp1ZxckW0mG8k68Dxx5MRk
1ri0i8ZsZD2CNbhebXhG6PqK8oEcIAdj6gWogBwDbDCgqyPoUJ+VFM0mY0zXy6iX
kQ2bwZQEaRsA3TcEmkVU+Mfxkd2JXGxkgH/5b6dfdjIcsML+6u0WTwXuMsifxImi
UaJoCh8682nZQ3BE7A7KIVmV2YTu0q+R6x+YpHx3bliw4TixZxXtYx3k51wtoZ9F
8QBcrTZvPbnMDhb3lK92M2MeuYnMDhOQULE3v4L2i04EHVH5Vb4royy1UboOzDoz
swWlq/8gG3PEe04Thn7+urQ2NRDjsVonD3hvQF8kfSrCz+pi0pccimaYmHY/rd/7
VPfoG1TL6FO0CwMJ+BXxK2rsDgMFZ6ZIa8WjKzKT0Z6qR34D6FK4G+xwghiEesQL
p7C4sdKR/ymH88eGvIcU/r4YZTuvNXMcBFaDKx6soQHnhhQwRvfFJx4JtGPBE+k6
oMEvY/XpsrSmSK1O/fAV673WgW3yY6QYGLxr1bxziqZiLKADZyG0F/DUfTnVXGRm
1iwa8SHk8azMEkDA9jRGKBlfk4R5tFXc+HgbIHbmiSMlSJShohHeYvuq2yuTy2md
mFCTSvnoUVDZGEjPgT75klb9MafGRToBE/QF0iyqHI9c+Hu8tQpVM5mAH3vdSw1K
vzo/7F2hQbvBYmsw+i+QZlNHPwGel7o0tvSxLjd+XYZUOEn5RyY3QL2hQoAV6QG7
Xk/m78It9EwGve141hFF7+eGV0Uqnkp3TVOyAs3zH5BwagJwf0lW861gNyfWbIQ+
ZKxK4icOoByMWo2PbGQJnzmdumoCsAi3YVHmmZpvRh+yQ3WdUBtvuarWIKStA6z7
tnN/eg9E5pJs+4jeDGahZrat9mMVig5eVzWfP0YbUqTNQFM7nzxuCfVxG7xe1sIv
YcJXco+qxpZlybdEjqSSN2uwqkMMuoCcxg0KX6FpkjhM6wMWj1BsQQJ8fEV01YYE
/CMW8rMzInE4+0CeS2GuErzGQPx8zCWNfZus3IKvZMlti9l1+UkhpywdKj75GpIl
2TBo+VIlxWmgBM49ySBM0ig6WSscVdXGHcqLzXdPJNg2JVDyZPIQiZpQ54jz5G/h
68zPjlwpyH3YND0NOPjYkcF4DjKKv/0u8t+7L07W1MiOqA+TYOTZMVoyUCfwgTNO
77FTqTbewHl1uq0+KhVpOIbYhNDxfuDe9vxuNIUmAlejqsE8hUG7TuN6BvGyq6y/
ckHcp6BqOECYzcX7HnoNhzLfs35jNsv+LF9QKhmJyaWzhm70SPCCFs3WeBof64N4
mOkm0NnM37B33RoaXElytNJzKbUSh+mSDtGj6p5z3i6044tbthRV1RkTz/HB2vwX
9AT+/yt0/4wNPNtbSXb8WLOKPhY0LsZwnWE/bxW6NZ8VJvUaOGnzUqxXgVFXLtqz
/W6hEvkYA7g8E0ZZTXEJkHZgEH3u46R2jIHV7VtxMOHRKGQQa5LyHIsVFMuvpPPD
3fK9aRE0a1lHM+f3pKDPBlMf41CIXd898AEeiS8zeAs+c15Y2ZMS93zMXl53MYYW
eb5fKk6znJWkeC692i7K0/tyhA3vVu7YuF37wV7JOkhpqej1DhutTBZNtXKIPZkA
M54BP9c9ABRFUwemxdFF9lYJ1j5Qvyi78Mh5WSZzRWB7aYVlL0rOkYR7t9riZEp/
9tro8Od2Y1zYKL2Od+7apUesdBBkURsyaoc2Sl2jSJS513Ip4tB2FmT4LoVxaWzQ
i1rO8BDEWVP9wWqJ8agHz2fYd/FETd93pQk/JUwS8uqEfwC0IFl5PUbGL/wX2cQf
7Al+V7QkTTkKvu/VcfVdthrTMrSrGHe3rDB089wD1lydjakqX4AxvlSG0VAFrNp9
ZWGClin7cK52X34hPFAPsySIkuncme5290aM5p2be2dUZqKjkavXFzADWSgbsX4V
BBo26xVNH4ZKVs1wtmBJplpEneqjjdrCVPwiDRF9TIMXYWoQjmNKIjuvVpqgM3qQ
b6X8EkE+lyj08ZJAY6hn/ARp8USAYLGVcmdn8HB5cpW0WWInbnYkzmktfVT9RCMV
wZWLlTz+jloGrq3KSeN1pMot1tC5/KK7IwHDLwfS3gftrjF/JAhaVyH6oFF1XIPW
HiQ933d0NwudIw4+uKK1duZu2g+3RYmRoFBUL8xCnTwrhQ9pVuelI2ISfIj76DQL
PJg2Xyfo08FKayiENhEiKI1kOyWeiXtVNqFIfRjlOdwieYdoutpnYvRu9+GcfNhe
HT7uTlNXV2LReYOWh9f00eO69ZfnazGA1Em65uSz16PEnGmYsDKczH2YOfHIR06a
E1GcB8ffjcxw0Aqxwr/e0/XM68K2n/4ZcjQ38KQWLRoP0ngbNbnSPdS1/CaKN7Zg
qGdWhWKJPHCHR8MXQm5ZPr/zIMt9/YERiEFXjSVFtqbS2gyhdei0PvCTg1CZHcTY
Gi8KohU9shaC4mxlZP3w40emcbS8k0pAcievhMH9FQqZeT5bUaxhZLCJuImtfMdC
TuhMuj4qEw2+2HQGvTeWwEQsilCzIKyVeSqbT3vDtgGRzi+ELGVoWQN3NA/yMr7d
8raBpduJ8z3jewePRyZmFD893GlVIbvMLSDUJG8GamwyY/yXqE2wFyDNZIZsnCZf
+DM2nBNkM+f7axcr36iWiES4Zbp3c4t3pPiaLo+8B94qRFxXf3KuA3BHI3+n4YEt
jKPx1pkYnFtDnh9TCvl4ZOSL1GVrxMUgeH9MD0YzYx6g4b99RV9aBvFvd6n/nRVR
j+tgeyJDBCzy+v6KYjZ5hTGbj/1/Vj6dF4EgSQF41CWsAB485f8DB4OYNLCf/+RM
O3QK6NmC4zzaoHkKq8XZgHCcVJD32UDBOCHDhjE/iqz8YL/C+BogLrIAcwiqYySN
+TPvYda0vrNtrBXrXl/GqWzlyaio+ei5n8G2emOpxyB2It0rBE/lipfcIxVrnuzI
hB7CHWgT/tp4RM8uN2HoAptqkWapU/DfB6EhPaLu1aO7fVmnhWmihYBDe5LreEVD
oTouQL9zjdUdk4WcgsFD0UsaAF2IGDviPLqlN6Oj+aI3gMeecuns0lBT5Ptukl5Y
c0TAwHpDBWE9m687Pmn4BKogVPAI0a+T4Rii4gC842Sa/f+0xLq55ekcgR7PhQcU
bGylqFfCW0ogEP7WCa3yhElW4FLD5SM7pdJ1lJ+9qdzCTZIXKKHwDJAqRuSMLG9h
ptqcdk5YHANhaMYk12ZgQIAQ6CoZVhG5rmgNUGJiYTUa2K81a0sTw2ptJ7Nbc4cO
vrSlP2nxaS6yUCY1i8A+shd0V/CEGXb1EZK28JFX3mBwKEGhPEiiFV/67gxsujez
zZugOSGmjH+76H89soI8WbfDBNxa3c6SNaCwy+Cb43ada030gvUzCYY9TisTK9B0
wy5Hu3lNntrj7w7+q3JQY6O/WvGEPT8wCsVO02DUP8c3/z4r+wq8XhuGd0Ex+TGQ
b61c13q+ysVRGgjWcIx4kJIl0dzWTmYAXQXC7mK5BN2rJC+KBKtWBFO4sTH8db4j
B3N9oZmZB+YmzayXapLEbuPEhCLOOQo0TeXyTfbQsGxalxgyZU7A/tUO32Z1gJ+V
rQ5avw+OMeS0FZGRbb+QtO1S54v0uoBtFdNvHPxH8+7L1bjHNrlJWpX1yhhQbttv
jFr3ohprKPBbhVKiuvyhwD1cl5x69yN0Pw3DYBMnDOdrBO0kEka6qDVmLfFZd0Wu
5BBr+MP/YrGsfvClfeWev+m9rRVvfwFQtgFPwIFeCFbmO6xnHV21G4cZ9wwPFzeI
8TEF8ynQle4VzTtVMxAWeRN4+9A4ijibZClxLOZ2IMFI9PFSl1bWJDLIKUy8ihAm
dy6gFbY07H4DqLZuniBm1+Ocidug16wb4XYrImL9H1NcryA5JSW3aEd1mRxhP6S3
NbYVFKFjDi1D7dMdAjvcD+mFA1pQffLq1Mlker4VhHNKk69L05p3vRErSwYOFvA8
3auSAkGz2+9xGFhIrJMwhjw9Cl6N64W5Hla8Hu5PRSGFabLDCmHjS4HDzZNTa72Y
njyreDr446XgJdcxiY2pSC3NktYXv3sI/07hZbPo/hXN7DHY9lmanGYex2pmPufE
0rAdoAQi4LVWubGQsbIe/htoiK4COhsJjzlotR2TYDS1OydW5M7nicseg1Fz6Io6
ixuxwV2H3R6lxdafvQmVms3kM+OMiiTi78xNIJecu4+YgIogkZoUohxWArSb5vLD
MjbslcdI1Wuccnz4m1SYPZZkJdicMArTFWAMqY0CYvYr4NrWdLzCLoQwQz1CMBdP
2X1GIC99PwY/HrDFH7J06y5+ThMRdUbpRPm443bN4TwVz5ctA68pH7R5Ssf5ZQj5
MzRa/+yzP+quj5vvLZKEEBN23wjxd2G6cjCKsL4KNAUBvAV3bPM96e6Yjwbuu2le
4smVPkELyx1I1jy6Alds950b7QVYsy0frSJTZJI/qVEOJuxyOdgTilLFgRE4eP5K
9IIcAao8akxonMvrQE/WCw86DlwGgOa4bqMPOPSRgk/8oBVOO3Qg8Q8wNPFhXdfy
Y0dOsr2WGjoRbAbeEJEvLLK0kC9C+xqmLvTe1BzkMQG4EUqSLn01N9KHdRu8AEW9
xA3sFnjOkVsscKSiEpk8HVGiTge7byJPWz76sAxA35EId+aDkN6QDQ9FuQgkYoXn
oKQwsfR3stLkIj3umJOAgCFpH87KFHysqyAm+7Bici5S3jR37IEk1w3dMqXBkJvv
1rI0xes7XLHkte2HOhLj4afqNNRELxbvxEriWkZjDU8GddfjLRnhplFETHBhqGt1
nptNKM1DNy+xYjycYSy1hdYpX+jSwYjdw7XfHTiTpaHxVFweQNaqp7MSog0sP+Vg
5qtcnVwxYMzANj3ylLHZKFQgFoGb/6wCGeBro5Qg1Y3VFIHs1oHzBM+ToPrBCtBZ
7FSNYY9KHL6SbC3QXz04gOfzWqLEHt7h7ejS1fqC/bOenLcKaPKGumKMd/BSnoCT
phdwGBPKf4m1cjqj8zHCzEls22J9lslUu/KQywn1nTTlhdA+Zu2jxWvEHLI1R4eD
FTW0Y/OkvXYAlnFuDNQN5w9kV9/XjlAbISf5CxIAGkbKOAUafNFFWyZBmbdaJ1aC
YVITEEnAXtpCRnFP0/rGQsw1TshLoTlMnja0Np2NxpBnyM0qnQan3f8ciugZSyg8
cHChhGM7vFr4Ryw0lAa6fOXE0vbHC/FAxvD4luZbR1+b0pWehd1ILhN+I81MYJjx
FlEkmZDkKZMguk1jANHgR48JN/dOZl1XMb80adKH0qZ1SF1ZD4pQPkclL1Wn0cNt
A6RdzFH3wHv0AFB3d8mT5equmkLFiLf7cb1HhSprbPfgedgv87ZrPGMAYiBz8lLz
ZQMM3XNLavRHQJAM+AqtxE92MqsKVRm0HSxysGALwZDJgiCxPV2H3Qr4IxXYj39n
M4RCxL/HmCdCM28wFYM1L5Z8d3Zw3oOCzT73qMZwVF0aFgjFemkhyMsBTsWWn/ls
jCtRdS1hNmd3/AWqX/Ec1W+zeagVw8QYiwdFmtS8dIEb4+2jq1tc6XNmO8Cx0jkR
UNu+A9WuOwWLwVCCYx7vX6IOH7U3gEQKEROJDwxWM0P4xuxObfuuIxPin6eMaNg1
ercB6Si2LzwhFlix1e5MdtRwfTWoadMLfipTyej0MZKMHj0eyTLwHJ5+LRZ7/+Gn
Al8bZ41c7M2uRZ613sXEb6s40gsrFrpizaFBDOk8pwOvg4lGSDOkyMeP/mVpXo/2
8x8FJZnSWYsDemDoOs8+SusKfJqQf/MjiIQBB3FFBJpYEeHYT7JfSlD5Q5RWKKJt
7sf5sCALAKSEqvM80sHS83k/v347iF6N1qk1fDU9UwemU8lkVdUPVg2XB4GO2lgx
VG8JTw/WPlOeSw2EsTGorv6yZV0fWtPkoJD8cSFIDMFgFOKLDkjJMUN6umDdD86n
PltWIr2bzeUNkv6utZG5S98EmXCLY7TsHy6/D49LREC+73uSWU1Z5hsydO8UEswe
p5sp88UU+EpUmFNqOehBGWj+M2HnmMi8pCqoMcQdq0L32YDG05dJUohL7WqoKuKK
dIX0CqWb7PXt5RVflifirHRw//4JkNkEVW/DPrk66cuCYrgA4uEewC4uGAzuRGpW
QbplX9tnPLVPex/O+RfH75cJvlEluB9Wm4HDjxGUz6tH+2if3/W70qhuaG1Tp85C
rckXbRd1yrXWtQTRcBl08XdxBEydT7IYX9d74/Yarpji8pbxeAix2MLO4s2zwPex
CbJjDi2/5t2eBKdfi65KQTVIAPXJyvLYUbCJaP/CYSTodEhEbJy8DHJPaVXSfHMZ
ejHkJ2GSbZTVhdpBGunpMnoi0zVXnN9tXXMwDBCRrSxjqyJvLWf7fMGNx0AYIuE0
8tx7rTA5ea15R+zNRMf9pnDQInZ6bGvCStVP8braa97h6f7dZcnzoHzljMDb0WzD
FP+udvy+2+n7gDiZ5DriK74hBmLkm+8ZloPorn5Mj+/AerXIX/dSSh8cbf8y7R5m
aFS8T5OCt0CUe9IX2XjUmZvzTKxW2AkF+D/pVG3ecANimWpY8iltJY7VNaMNkiMb
Fnz9rLDPWNqc43mGFUhIwnj5kM9+CH3XVMfYuu+IvMOm+sd8LBR3t01TDglO0iw0
z9ztKyORHrphY4Du+zcUys99zPkBA0A15JMgyrbK6syapVl9E3NLavuhFd4d/7N6
poLbLIdwsNixvXrh1nPcTEcETVZyjqZ21CmG4bwiFFbXYJG7UAEiH3OhWmEKaoWn
i4or2ckcG1tzsoFZGgzI1JfceBDWDT+pC1Fer4nIjrf+B3+04LLE5KXI+R1XQowl
OYAW9LYEa7bvs3U0ehFgDiWjSrEWttD99y6Fo2qHIS+JRXLSakBukfKIRYnWqtKA
9ieXwFd9uVbGrI2rn0jLpxvT+Y6RnSsJKL7lCA7OzN1FVkEpmTt2IfKmXvxAarRu
3EpEVODHIRfY2LFsAVAXcXufFeO20nwdeJMOHEJStztZN115hPOmPb5veQGrTgyv
tlhTbDrPMtDXPdxnvmw1EqEljNcdaZaudP221DXnXqgop32uYL7QUNfxFNRo1SP4
C0YtDjsBACFkaq8zEyFEFC1q+wEei+gt4xxdq+Jyl/8f2gkgkVbSpe9DlYnr7sFk
lU6UPMfkGupXoZqUXixXvAmuT88dVwRAvooRbPEQfNHZm//shFFP4jtFFqwH1Zvp
wJ4pyu7/n2KGTMKtewanC8yJFzY0M8nsFzdfcNuEBRk1FMxX5CLygfYBzEuFuXkY
8Udjt0Z+2TzVdMG7zKJIiWXz2jVEwY4LuwZZmp/2jmmp4EyAi8hkaPKslQh6CLLD
Grhc/yHRFO1RPra0YTogDjtfLt9ZeX2qcSQ0GYmscXdDdrovw4/ZvcxCHltmdjl0
+AoJ6Dtzc9A6LH0FKG4hqjVKGcvrjVnXt0hY1b++yrJ/WfrJvs9rAYMbOEGzIEzU
P8PZNeC9cEC0kPthmJqaYb2DXP6iEVI7d6qzRJzF0kOKqHHlbljNITSFmYSHapyW
vNan79/x0/4PQM8T0X1vM8o0zBb9ZJUOubehe3Cgf6N66acuuEtWITOvzmsP+F67
XHONoX0GPXnQoOJhkWEI+OjuxgI6HjnU0r/zdar4khxNuovlMfO2LuB5wv3WdaIm
zIdIVrJXQASwvVB7347JS+a82OnKINJGvy1Keo+nsfpVlaO9nvJ6tLXUdA/oEF90
TMgG1s7tpayAWEIbOoLFu8cB09iU7imAEv4d88FFCNOCJEGwp/B6e3cmuR0sRSRQ
9ecyclebpIM6dluvzKjWYUTw6Uift9GPiDonlP3Zhb9z0ImD4uH8KDyb8ROPCOYl
eaydx7cggJf+VODJ03cgfdo6aVPGqxjG5mIG+ua3d5Bf8UM1Um0q2sfZ1lERjcaO
e8cMOj5n8kMnUC8bdvYeeYID6wUrpUEL4hCMKw6Q0ntPux33cgtsochAeaWBAmDh
rem/C6wAgypQ93V6F/IOq6Bs0Ow7Tq9B0zixocP+GcYeGqbl5Z8xNTPA64DviJ3t
mAZ7zef+naXO5bFrgG/0JVGGF3w4cuqarN2B6NqwaM96a5kKkQAoRF5wdp7I3kZ7
ggkBV3P6sRWEgpJaBFSQOgd5I2JuxE8Nezc4A4WELF/MH1lHPmicg7amZDcBicAc
LfDcD+d9v9wUR7CNQkg8dk9wYQeIasw1MjxvGto93f7b0uSmA6mEQocHIdWdjuA/
OuSXlay9wzu+kaAGfu/l47bLR1QHsY0uF9A8+yQ23etDECqn9UXOzJbw++/2HB3E
+/m0sznHRDB8HMo5jbThve0hOXFS980wCeDCT3H55jQliKlDjbzpHJ6mlYmxl0a5
YZp0squ65MSjF3KjH9qpfh/TemCc3ZGyxrQC5rTbpq8smBGGJ6kG+2QZBCKxm6Y7
fvtiEGsIQ5jWpCFP/m60cJxGg7i7M0qsVwiI3vszXpUCOwsw2pn5qTw2NLMD6OGR
d9khxG2wUA7m8YPV/xfXSQ4dCQK6eW6zN8xNG6AwFNlldqhApNNn3N+x0GBV//Mt
7he16TfcQJeyU0/YfpiumoS0pdB69IWyOF9I03NXozfGLDvQCc5ul3O12CRAGfuD
kn9ZtHugLugT9pTVKPNw7ld3UbTUvvRIgysLT0JhAFjEpCao5KIkZhTokVQkDLxB
jcmdyKnokyZ1kGnfJ0imtKV6NAYDi7MDrfmvuzfy5sXe0oTesyJMGipBuGi4Q5C9
YJS9gVl8GOSyrLrbE5IChV3MSWcAMSaMxd54fJM24+guteT9q/xOWliI8BbJqG2d
cjqLUSWw9gnL4y/dpWV+MelxwFZpz4L7OCV90FCnN0jRVf7IQrO0aqFlg8zoAgLn
eKWOPfY2Q51REmyVQZk+ZTiZ0nRimhyU0FsTTpaG2odiXmyMK8grwym6fRmtsfaa
2olyNkRVDyXx0yIYs5GkYYcYEEYuOhOhgHZHKJV7OOGFrrB33JSwnNkOhy8y491i
Sp1RQMwp4wVAp6OdRwwKl3ijlWX7IgJ8upEBL/w5+AfsV35+oda5NDRt+dg5n9TF
OLbte2/gfKGVnQSxMWhgWC+pCNzfiuHfvwAqcBHARcTN189YAPYamXxFiojvmFvu
QBwXj/H41dfqAowNtC4vhpe53Z3YPT0jbA6lvJX0IgJ0XgsibBCJMFxj7oeUF926
kd/mWA9Df4JEM+RV0USvm8mz2MCYdXQLr4o8BJXN+LC9NFses0W9/XOFbAXT/gvD
/38ErrdoZCNvhtCkqxMKrJJB3IEQ3CB0ezd7esSx94FysPsAiPzPzIDIdwc5ALJE
axf4UVMgAw0D6Gllj7CcA/Yuy8NWoqFlys2P2kOFBl+Lm/lP4QUTgKWw/FPxX/4h
0bwW6elux55YvMKoibbVAZs0BUcSqvexW6RZA6FSvg6zxUoNLcYoaM9g0lTsmHlr
is073Ld4XR3VM+MfciiFXjhb60UDcBem+Nqt9hAf68r372wugDZ5TmvdCIPwhTly
FJqMrzItRHA2afoA7i/ru5gJ23+DCxVRjV1CkqZBA+WKyAhzp21rp3t2GFFJPJN0
w3rrds7gcL+BgDqkF4EGFp8WujxOwjuX9qkdtS9rrXBU2JDHat7tIo3frqX9qKqX
4zlLOKa//3X8/sVSDRaatLETrl52lTTOd3ew2iiqhq1vZcGGSndZvw0qhuzZbWV5
ICH8d6JyvCHcm0Nos8qp43d6/R/d6UCH1MBcVbopahFUL2o0IRzSxX2JKIlX4k3G
7u+i60yfIqzYt8+Wl6WWWFvaYEMcUzZ2xx2Icyi37Bwn4npQG972pWfRm6nvR3p9
iRgYNGZR1Z+7kY4TEZiIV1QEDIba0PRM+GBtKxDCND2DFnl0c/FcjljA2RPvqIOu
9OJs3dV7J0GETB/cGO+nI64onUSQZGxLyn1UoZO+OZQESze6Yx5MjSftj7akJHGD
vJL0BsD5t+83OozQ3k7DjKXF966B++XGKOCCNVp0Yj1GaqRwqeKFySvPGIWPKVvZ
zo+t6K3gMuFm/4aX5ud4amy9ZmrjLXNzyLYKHSHLWLREROBQiCCKqLJghODIYBzC
D2lMStlEwjPvbWBlMpD+EUFotGUqd9/vB7D+pYX+60yL7SAb2WaJV+Z7d9CB7jEs
RU+DOspopYT1lFHCyPP80ePKt8aNYcJoOVIBdYu3bphtMPftYfFu1ZT1S1upVoCc
8g/LyQqmvmmpdwdAVXBLcTebOLaPtYhHSqhOuJM4VlBllFBGezk9DWtua8huELTM
d1oF4vItBm6YQDt5ygBxF2XpFO50RutDku0cDtq9nnll3sjKUw+eKEjXjN6j2PYk
+iJpL6C/G2CLv59BzsccVcdUv/cRtWbTf6sn+maXzrOKf7en3PXGxK9q5YODHyFi
B6ILjo6YLQuR+/EZ5FT17LO8JmWM+LeVIc3CkHa53KvajqhON/jybh1FyUbT777O
O7Hoyh7TALuY+IDRPakP7zasWzKnuSYVHDZTFBTlINS0bIv4KGnXq4bY7vt3n189
7Mdqpw4Cbb6lsnemsslaZX+Da10LF93g90PKl2CbB5Xjd3owLHs+PCL0TOjmycW9
8EOExhROS72JInc8jn7Gux64tmQnf8krrE9svl7Fnc+VRH7+D9UiU4Ea7AYlhNiZ
kod/3Feb+42cuWhRw3mYsH2a5ncFCopZjXbrt6f+bT3LPERn5Fo1I0PaVm36DCto
0R7ye+EtP1U8os6HvopRPC9zsLlIBCGic0h+yHGRtCPqlCK0Ct4UYCVJ5KQLelS5
LLMbfCoyhE7CU3wOb2nX8U2GqgOIrXMp0s5PVqyz7jwmxylORWhl8Lv24OCYzxK2
fZc8OdYrdX3r+CZG1q484RG851inSIiw49PhGkefynPYvakc59RPJtJSEwxZbJY9
+Itvjqsgx4gG3Y/igUYp/gtxpeGNWAuHe4XHzSHK3vY8Wu5rnyHzmXWvNDOsby90
TZhcPLO/Rv+y5jk4KzGVQ5p7fMqtIVpb+1X/+iR1ddiG9cMIG3R3Ol1FkT+3McYF
DtyDrXoo2A9pLOA/XvK7b0S8fjv3INjM4Hn2tIvMRVkDHPp441qmMMjDgKs7CfdN
sfGK4LLy197VDuI33Vkl2iS4pxEvWkNGVpHKf+JZbp6AOsQibIENmBGsfviw/HP/
9Z2UPDtcorfWumHydYPPEA+JIYJEAnn27wupEV4qjLrKPrZ7btoUKCvcFiI3E7iE
xdlTngKs5K+wbgxvHSWjhLVQbjvLyLBmmbm0ndagnd2XmUbj7DYrZqaOrrWquwzX
spwfhKwqKUSOBbmcG1KbE2UrFabvT3Hc/YNhzpjLB29yi+Sno5tfmDmmz/ellcvE
GRjPz/1kLdevMRVaJ9ZC7vPFzAuGslS5ogMN9LUDqswff6v9Fg9j2N+Xi4tSAwMm
EmWyenqxCJljpSQeO0vw3FMtgtdTaNsXq8V7Nc7ds9hU0hLDmlsLeaf1Aqz6DdFr
AUl+3m/sWeNnPaE3ImwsXBdow5x4Y2F5fd+YcR1paahcxd0IDyZiMhe+QHn5BJta
6R5terbSMQekbbBlAFoy3bYC/b+W+Zk4LUIOqA3oE6FYSmI7kqmk6DmZHgL3TD2U
6MYxTry2oqTEawZe/dOjplFNeSp+twTNi8Chsv7lYE+orDfvH3BQ/SLMMRFi0utr
Bd+U99IP1jSF7VeX4vscdQ5q7j7s7KAMfvDn/4vDFXXJ6w/ka7J4WeFf+xvVQCqU
mLSiBp0KtsPD1QU7w+jjk2NCESLpapPBWPyMaMIGzypYRfM+DY7LEcCTJv+xmqAE
IuqsBrlEgmQnm7IGyPg7MVkE8BcRBhUjlnD+qyKSF8wn0kA+jy0XW15tIBsx6Z6G
y2J8AA6JXD17ep6zex+vqK6ZAGwTFCBIg4KJ2AOWELDZrJB+bo1qOHG/IyClqlw3
WDKN4E2ygxd12Tlr2KJTgXNYZrTpJSmyU0XB66mS7LXnsiRMZnaMFI+XMrN38CME
IJKDjZG+uzOIOfZ4kKftrckCAVM1HJ0F/i3zvsuJjjY5MSSGryn1umWJ/ICbpL4I
MFq4UtmzP9fxWWFcQyOHyawQdLjv8+p1WdjYurDe1kDlCQ94BW9cQ+HnTJT/7iK6
Wj5KHJOpoCDmFllUmTFSsyrE1sZujppyNxotcCLpjCt84C+heYscMJEi8ssECuIu
DKdOtZ8XeZKtMeY1o/ozPZlCRk+O2qb1WRnt40SMffImfwM5GkbpVqQjRAbQzk5v
QSGXvwu4vsjchqp3lRoS6mWfcJnimmdHOuTOdJ6vtMIUU7kQ3Whe4wFLb3jALzm/
v9FJJ8bIeGVpTC48J72tAlPXBeAviFJRY/qK7WswPPxZrCZGtY1opEA7eedrIB1V
QkS9MZ4BJwNTywVY3is74QYwV+/CAI0NpOBuM8bYXHLMn5jg8rS4sQG4HFnQJY5k
UstjIluzl9xI6PbJmEl5kHFuFsP5KSH7gPT1ht/ssh/TKzRheaTsRN4vgMAn1wBz
XIjCO/zQfF3gNvJI3SfyjWh0L6RgxC+czk8Uf9ZS14c04JVPE7hSylHwzL84LZ99
hOmFaE//9SJS6wflrb5O+nAHKcwpeu+k57ska02BC/wKpJFEAJ3FXDiMxSX2Qhl3
u78GcnUvqagEz4KWxsgIleLZKS11crNcP60U0RbGmAAQNdyiMPwkxJFkIg7D6cFo
5nHPci3gqCNm7lqC8KX/aNCd4R2HrCCeXM38gk76H517oC84VvxFzjNo6/u8sGtD
HZVQuA3gfHevYbzHTpWrCycWeB1EgebnOuEg3ZhHmmad23U9iM+Vn2Dv1kPAh9zL
P1EXw5Zg8H21xTQcnBsroOqz9P/ZvEJ5ClC3X9vfx0SsgKQ7aPrXQSPOliGPj791
cpoGv4hju317ALkdXHCRe01xZvE29WXp8jBCic3a6DsO4MurT0WtZPrpMj04DYAx
fPecE8j7ne17Zv2FLwFsIWjNVz1ajxm+VVQyU6DmbAg3wtHrCoIN6/t8zPsvxUyn
EM0ntwx0XbtAOUriEFBN06GA2aHMY3COJEqokVw6jo7V5s4dbNW3x7I7M4tU2R49
v6GvuA6EXisuiBzFsgFf+MGrZlaqFkGIO1THrjgLudgTZXPcO4JhOK5LfmodjFSp
CnHcUf8MUE1JMTw6PkN+m1jRPDGrLOcMdEKudG6uTrIR3OyF9/j6dibUk18opbyv
ImEGjoSropLN0AgN/oQa+XTEWXrPt9LyUosQu9L5d3nlZfsbwmwzYPUpCJP43bDm
wWXT3MHujTml2B0bjvGKJo5a9BYbwojbH5eqdBf5/QvK0/KIEDn81XFZO7VJ/8/h
bDTwLCCnynFYLr2zuT/60ZcaH+qGVvntfH7TAc0g2BQbPT0hDmtSSpZQ2OiqXdN2
rrmcxUASuJSrk0eb7HhE0L4fySc/Q5Q+56RCCakCQcH5fE5Aiez4hOjWutsJ2BA+
vtqUUq/sWzIWQkYis8gbAKGvpMzoYSi+ri2aZlrXxYreRBOkL+HAO4X4/5dEBwxI
fCsSpyWSgb/+Qd83oFHCg9X5pCnFb+5vbDzgtabCj7vNLuPAeuTbz67RHTTbcX2k
9pOxUvHcQEe/GpOy7mGenT9LxRso3aKvINKJbAqSR89lbLnflVOqFIuUm9/ggMSO
v7eY9L12qYv8ZQXQlaNOaR3mvIAsScDlHEcOTRkqQX6U4CXorrOJIOvJmYFw4QW0
kuvVSQz69Vi17UApqKs2/fnToCevhU611iVOhcuV/Hg1Qmwfodujfnod4laU8brf
eG8lZHnDud+8ajaf3BQ0uhTXcZvy71zhmHesbu4gLQPX2kqE2Fci3KUvvj6pTCEM
n694nNY8yM/3zzhSxKWZVuBuLW9HtshxP2nUVzNFcbxSCPwzJdfiXzKauyswyPVT
Qrb93csSLO3GWzBP/MF37Updl0oLW6Fu3eZf2BpzxGXeyWNOrGSfxUwjJ//uWmtg
/MynsqQAj/DXvXlZNO6olx9zWkCyLaYz+pRCkEVOeqgWjc3GXEtjYPgJ+QRNaEDB
R6AmVXv0ZCO3JuCzQXVyKUOc0KlSu49AbgqrDoX3606A9/HfVsV5GQyQ+SJ29eap
MJG4czDM+71N8KCfNQz/lXt6s+Jfu3q+ftIOrxyPyTf/7isRWPvYia7CJpqVC4TC
f5vONbh/SVKGAWZieX4sAqW8kuhtkXretnhlaM7jjtA0HynQ18sSu+mRW4RNsX75
8TPP3Ebkle8xvUjcEpDuAngIpoYKPu79lJ1BK2nFzo07ZCPfLstBfzxnlKUnlkQD
UHd1YgDvWPTxr+z2iIs6rVML4rhdH2CppK/78d6IZ+Iopeje42mVMqQFqHCcycic
n5iLOV5Q1sh/Lpx78YR/Lg2rhdsGbGQhQr7MVaG5IpBk0IBqxLLJ5w8uYKjve4S9
aoN5Cp/Xjr7iAXEyXEfJ5Ww0SqZwNLb2HirGKLHQ/zHxlYPs35FEMM4v/SNlWDDb
QQTpXw9QLzfCW02oarQ63nnqjO6qXpmX04n9ZPt/FTMZSwrs3Eedc0qyyKTPjH28
JHrHfsHco+0Tkpm69HGAOBXyv28+edkiNYWxIrf8b+Du3ltwNbUoiG5WqpWolrIU
kG0OhNsC5g1noqtBdDRrCBfEQNiJqCdifu9MyRClWXQ5MAIpp7IohHnuFp0zaHL/
kg8lP8BRKaoOxOgjrKMX2BqXPdywaYuNZuGFBHW31Pcu5+ySKTPO6ACWyTTGBwps
mvxTvxpdQJz4Mes3xoVJe1U9M17lfJCP2ijThNcmD6r1ybZoHoiKWoXCuZ13K0Ha
y0Kl3E3D/ni7lxzWXYj/3pxR7C9oit8eoA1dP1c2a13yA4wlpPXowrflntpGehAQ
SyHvOCwTRdeFZzwTeQeyuNuQYY3ARyfh3LxqQCz24L4SNWa94NKuRAUn2iz/L17I
OhGheC89gXVNKFTjlbaHG2lHeCCv4F2cryowpa5EfFyIibxzkLQQKY5Q3vwhCtva
cPDxc8QYZlDTAoKEbz+fMtgfuYCbCZlcStUqVcF5qg36nOrHGB5/lN9COEn2hCft
Ao4JiqokY7eqMSE2DWIxWMYVkW+8iH1V999y+FY4p6iWYMbtQ6Q+LAM5J0ogyoah
S/ChoJM28Yn9qJK6wqgcwmZ57gdJoD1f+TDksy+RiKbv7eiRkBsMcbcPsUGVUQXS
jNWYessb7BLEFJyyrGMmjApiG6Q0CCev0YJYtzHDa0QTuBpLxzY7n257QQkU4qFB
SZg7PhLNxvjO1Fbb0sRxEU8EB8Us4UD3VX8qY++U0T3DvRs2vWkfarxBOhbc2nc1
chK3leV4RNVVbvQZHNZ91aTu5sXunRfEIy1XlgO+ZgY/1aIV2kTz3Vf9WJnEnJkK
G6MPRiefGeIsz3bwovOhlDuJLcWjtWKItYAI5iUcS5WSDoJpZaf3+hdOqEKWFCqd
jCHCBIpx0JGHP/Xbo30vGwxcDzpOOv0tYWmLp+CrQKCF+VVGUO5AsFcS49xdKCew
K3Z6CBiXvBjkdlGA9r+KZ/ZXtvZYYsdWJYLGGDt05T9E1A++vArAILOHPD1WQ75K
RUvFMK5pt4dcCP8SEwuc/gXpkVTwYh/ql1+v0JE66Rk+Y6bUIYlJOUl6BKu8L0qW
1J8vFjZ0GDA/SJeQOZEl26651x407hKcg4kMDQ841q/mUVyYfQcqITXnIDcpksDm
+uCF2fIZ2g5r0S6l5tLZu8BgAvNUitKftiiVRIeH+dL0mo2KCtIwxAtg/Jo0WQt4
0EHQG0ifh0vZvm1emLTRtIF1WMZUWo/tZRr2R4pgE9GlCbg4VAwLKadLNFF6vphQ
zduSs/5Fr/gk09yZibygs/px6NPW9a5d/TTLsP7Hn3ydtC0ZH7tQdWTc/NNg6Oew
r5UcfoYp/YP7vfWm4X3NLyD1f5RpiSyiLI++vql8SUO6fUksMZ/qAocZbhcRrKoQ
6Gk3MTN0Qny+TSvmOsv0s8dDO3+vW16Fy3pOHUqa5+hR6bEuXUKf4NPwe18e9qeH
LxFPB8wf7//EgVdgRxmomxddGwnbcn14xp37l0thkuuZUIZ2Sok/yW05ok9YgwKR
wCTCE2WYfvwiMkEfWHw+SNU3muBhifyYcuzzZMSHqRvFL/aqYMiR0DxCfFexfdAB
oml9ISerVhUPCarrzs3SWVoehHT40FF+Sqdvg35ZuFo=
//pragma protect end_data_block
//pragma protect digest_block
zX7tp1LN38+seoN2R4WHr/f2vwM=
//pragma protect end_digest_block
//pragma protect end_protected


