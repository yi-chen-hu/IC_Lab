`include "Usertype_OS.sv"

program automatic PATTERN_OS(input clk, INF.PATTERN_OS inf);
import usertype::*;

endprogram